-----------------Laboratorio Digital------------------------------------------
-- Arquivo   : rom_angulos_128x24.vhd
-- Projeto   : Sagarana
------------------------------------------------------------------------------
-- Descricao : 
--             memoria rom 128x24 (descricao comportamental)
--             conteudo com 128 posicoes angulares predefinidos
--             baseada na memoria rom 8x24 descrita pela professor Midorikawa
------------------------------------------------------------------------------
-- Revisoes  :
--     Data        Versao  Autor             Descricao
--     24/11/2022  1.0     Bancada A6        
------------------------------------------------------------------------------
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_angulos_128x24 is
    port (
        endereco : in  std_logic_vector(6 downto 0);
        saida    : out std_logic_vector(23 downto 0)
    ); 
end entity;

architecture rom_arch of rom_angulos_128x24 is
    type memoria_128x24 is array (integer range 0 to 127) of std_logic_vector(23 downto 0);
    constant tabela_angulos: memoria_128x24 := (
		  x"303230",
		  x"303231",
		  x"303232",
		  x"303233",
		  x"303234",
		  x"303235",
		  x"303236",
		  x"303237",
		  x"303238",
		  x"303239",
		  x"303331",
		  x"303332",
		  x"303333",
		  x"303334",
		  x"303335",
		  x"303336",
		  x"303337",
		  x"303338",
		  x"303339",
		  x"303431",
		  x"303432",
		  x"303434",
		  x"303435",
		  x"303436",
		  x"303437",
		  x"303438",
		  x"303439",
		  x"303531",
		  x"303532",
		  x"303533",
		  x"303534",
		  x"303535",
		  x"303536",
		  x"303537",
		  x"303538",
		  x"303539",
		  x"303631",
		  x"303632",
		  x"303633",
		  x"303634",
		  x"303635",
		  x"303636",
		  x"303637",
		  x"303638",
		  x"303639",
		  x"303731",
		  x"303732",
		  x"303733",
		  x"303734",
		  x"303735",
		  x"303736",
		  x"303737",
		  x"303738",
		  x"303739",
		  x"303831",
		  x"303832",
		  x"303833",
		  x"303834",
		  x"303835",
		  x"303836",
		  x"303837",
		  x"303838",
		  x"303839",
		  x"303931",
		  x"303932",
		  x"303933",
		  x"303934",
		  x"303935",
		  x"303936",
		  x"303937",
		  x"303938",
		  x"303939",
		  x"313031",
		  x"313032",
		  x"313033",
		  x"313034",
		  x"313035",
		  x"313036",
		  x"313037",
		  x"313038",
		  x"313139",
		  x"313131",
		  x"313132",
		  x"313133",
		  x"313134",
		  x"313135",
		  x"313136",
		  x"313137",
		  x"313138",
		  x"313139",
		  x"313231",
		  x"313232",
		  x"313233",
		  x"313234",
		  x"313235",
		  x"313236",
		  x"313237",
		  x"313238",
		  x"313239",
		  x"313330",
		  x"313331",
		  x"313332",
		  x"313333",
		  x"313334",
		  x"313335",
		  x"313336",
		  x"313337",
		  x"313338",
		  x"313339",
		  x"313431",
		  x"313432",
		  x"313433",
		  x"313434",
		  x"313435",
		  x"313436",
		  x"313437",
		  x"313438",
		  x"313439",
		  x"313531",
		  x"313532",
		  x"313533",
		  x"313534",
		  x"313535",
		  x"313536",
		  x"313537",
		  x"313538",
		  x"313539",
        x"313630"  
    );
begin

    saida <= tabela_angulos(to_integer(unsigned(endereco)));

end architecture rom_arch;
